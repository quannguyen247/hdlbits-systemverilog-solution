module top_module( output logic one );

    assign one = 1'b1;
    
endmodule
